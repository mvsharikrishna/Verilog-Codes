module basic_gates_switch(input a_in,
                         input b_in,
                         output not_out,
                         output buf_out,
                         output and_out,
                         output or_out,
                         output nand_out,
                         output nor_out,
                         output xor_out,
                         output xnor_out);
  reg 
